module general

pub enum PackageManagers {
	npm
	yarn
	pnpm
	bun
}
